module Control (
		input clk,
		input opcode,
		output RegDst,
		output Branch,
		output Memread,
		output MemtoReg,
		output ALUOp,
		output MemWrite,
		output ALUSrc,
		output RegWrite
);

	always @(posedge clk) begin
		
	end

endmodule