module tinyCPU(
	input clk,
	input a,
	output b
);

	assign b = a;

endmodule
