module ALUControl (
		input[5:0] funct,
		output wire[1:0] ALUOp,
);
	//为R型指令生成ALUOp
	

endmodule