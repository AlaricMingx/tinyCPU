module tinyCPU();

endmodule
